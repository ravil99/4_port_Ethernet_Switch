function logic [13:0] hash_14(input logic [13:0] bit_14, input logic [7:0] data);    //Регистр input logic нужно будет иницаилизировать
    bit [7:0] d;
    bit [13:0] c;
    bit [13:0] new_key;
begin
    for (int j=0;j<8;j++)
     d[j] = data[7-j];
    	
    c = bit_14;

    new_key[0]    = d[6] ^ d[4] ^ d[3] ^ d[0] ^ c[0] ^ c[3] ^ c[4] ^ c[6]^ c[13];
    new_key[1]    = d[7] ^ d[5] ^ d[4] ^ d[1] ^ c[1] ^ c[4] ^ c[5] ^ c[7]^ c[13];
    new_key[2]    = d[6] ^ d[5] ^ d[2] ^ c[2] ^ c[5] ^ c[6] ^ c[9] ^ c[10];
    new_key[3]    = d[7] ^ d[6] ^ d[3] ^ c[3] ^ c[6] ^ c[7] ^ c[13];
    new_key[4]    = d[7] ^ d[6] ^ d[3] ^ d[0] ^ c[0] ^ c[3] ^ c[6] ^ c[7];
    new_key[5]    = d[7] ^ d[6] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[3] ^ c[6] ^ c[7];
    new_key[6]    = d[7] ^ d[4] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[4] ^ c[7] ^ c[11];
    new_key[7]    = d[5] ^ d[3] ^ d[2] ^ c[2] ^ c[3] ^ c[5] ^ c[12];
    new_key[8]    = d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[0] ^ c[4] ^ c[8] ^ c[9] ^ c[11] ^ c[12];
    new_key[9]    = d[5] ^ d[2] ^ d[0] ^ c[1] ^ c[5] ^ c[10] ^ c[13];
    new_key[10] = d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[10];
    new_key[11] = d[7] ^ d[6] ^ d[5] ^ d[1] ^ d[0] ^ c[1] ^ c[3] ^ c[8] ^ c[10] ^ c[13];
    new_key[12] = d[6] ^ d[4] ^ d[2] ^ d[0] ^ c[2] ^ c[5] ^ c[6] ^ c[10] ^ c[11];
    new_key[13] = d[5] ^ d[3] ^ d[1] ^ d[0] ^ c[1] ^ c[7] ^ c[9] ;
    hash_14 = new_key;
end
endfunction


function integer eth_crc32_8d(input integer crc32, input logic [7:0] data);
    	bit [ 7:0] d;
	bit [31:0] c;
	bit [31:0] newcrc;
	begin
		for (int i=0;i<8;i++) d[i] = data[7-i];         //Разворот данных

            c = crc32;                                      //Каждый такт значение crc32 будет равно предыдущему выходу функции
            newcrc[0] = d[6] ^ d[0] ^ c[24] ^ c[30];
            newcrc[1] = d[7] ^ d[6] ^ d[1] ^ d[0] ^ c[24] ^ c[25] ^ c[30] ^ c[31];
            newcrc[2] = d[7] ^ d[6] ^ d[2] ^ d[1] ^ d[0] ^ c[24] ^ c[25] ^ c[26] ^ c[30] ^ c[31];
            newcrc[3] = d[7] ^ d[3] ^ d[2] ^ d[1] ^ c[25] ^ c[26] ^ c[27] ^ c[31];
            newcrc[4] = d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[0] ^ c[24] ^ c[26] ^ c[27] ^ c[28] ^ c[30];
            newcrc[5] = d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[24] ^ c[25] ^ c[27] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
            newcrc[6] = d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ c[25] ^ c[26] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
            newcrc[7] = d[7] ^ d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[24] ^ c[26] ^ c[27] ^ c[29] ^ c[31];
            newcrc[8] = d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[24] ^ c[25] ^ c[27] ^ c[28];
            newcrc[9] = d[5] ^ d[4] ^ d[2] ^ d[1] ^ c[1] ^ c[25] ^ c[26] ^ c[28] ^ c[29];
            newcrc[10] = d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[2] ^ c[24] ^ c[26] ^ c[27] ^ c[29];
            newcrc[11] = d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[3] ^ c[24] ^ c[25] ^ c[27] ^ c[28];
            newcrc[12] = d[6] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[4] ^ c[24] ^ c[25] ^ c[26] ^ c[28] ^ c[29] ^ c[30];
            newcrc[13] = d[7] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ c[5] ^ c[25] ^ c[26] ^ c[27] ^ c[29] ^ c[30] ^ c[31];
            newcrc[14] = d[7] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ c[6] ^ c[26] ^ c[27] ^ c[28] ^ c[30] ^ c[31];
            newcrc[15] = d[7] ^ d[5] ^ d[4] ^ d[3] ^ c[7] ^ c[27] ^ c[28] ^ c[29] ^ c[31];
            newcrc[16] = d[5] ^ d[4] ^ d[0] ^ c[8] ^ c[24] ^ c[28] ^ c[29];
            newcrc[17] = d[6] ^ d[5] ^ d[1] ^ c[9] ^ c[25] ^ c[29] ^ c[30];
            newcrc[18] = d[7] ^ d[6] ^ d[2] ^ c[10] ^ c[26] ^ c[30] ^ c[31];
            newcrc[19] = d[7] ^ d[3] ^ c[11] ^ c[27] ^ c[31];
            newcrc[20] = d[4] ^ c[12] ^ c[28];
            newcrc[21] = d[5] ^ c[13] ^ c[29];
            newcrc[22] = d[0] ^ c[14] ^ c[24];
            newcrc[23] = d[6] ^ d[1] ^ d[0] ^ c[15] ^ c[24] ^ c[25] ^ c[30];
            newcrc[24] = d[7] ^ d[2] ^ d[1] ^ c[16] ^ c[25] ^ c[26] ^ c[31];
            newcrc[25] = d[3] ^ d[2] ^ c[17] ^ c[26] ^ c[27];
            newcrc[26] = d[6] ^ d[4] ^ d[3] ^ d[0] ^ c[18] ^ c[24] ^ c[27] ^ c[28] ^ c[30];
            newcrc[27] = d[7] ^ d[5] ^ d[4] ^ d[1] ^ c[19] ^ c[25] ^ c[28] ^ c[29] ^ c[31];
            newcrc[28] = d[6] ^ d[5] ^ d[2] ^ c[20] ^ c[26] ^ c[29] ^ c[30];
            newcrc[29] = d[7] ^ d[6] ^ d[3] ^ c[21] ^ c[27] ^ c[30] ^ c[31];
            newcrc[30] = d[7] ^ d[4] ^ c[22] ^ c[28] ^ c[31];
            newcrc[31] = d[5] ^ c[23] ^ c[29];
            eth_crc32_8d = newcrc;
        end
    endfunction